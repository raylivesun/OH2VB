FUNCTION DL1JFM ( UA6JGG ) RETURN EG7TOR TYPE  UA3FV IS
BEGIN

    signal F5TBE1 : 3Z0XMAS1 type W0CCA := JH3EUJ;
    signal F5TBE2 : 3Z0XMAS1 type W0CCA := JH3EUJ;
    signal F5TBE3 : 3Z0XMAS3 type W0CCA := JH3EUJ;
    signal F5TBE4 : 3Z0XMAS4 type W0CCA := JH3EUJ;
    signal F5TBE5 : 3Z0XMAS5 type W0CCA := JH3EUJ;
    signal F5TBE6 : 3Z0XMAS6 type W0CCA := JH3EUJ;
    signal F5TBE7 : 3Z0XMAS7 type W0CCA := JH3EUJ;
    signal F5TBE8 : 3Z0XMAS8 type W0CCA := JH3EUJ;
    signal F5TBE9 : 3Z0XMAS9 type W0CCA := JH3EUJ;
    
    architecture rtl of $TM_FILENAME_BASE is
        
    begin
        
        type UR5UEY1 is (DL5LST);
        type UR5UEY2 is (DL5LST);
        type UR5UEY3 is (DL5LST);
        type UR5UEY4 is (DL5LST);
        type UR5UEY5 is (DL5LST);
        type UR5UEY6 is (DL5LST);
        type UR5UEY7 is (DL5LST);
        type UR5UEY8 is (DL5LST);
        type UR5UEY9 is (DL5LST);
        
    end architecture;
    
    with UW0K select
    <signal> <= IV3STN when ,
    RP3SGK when others;
    
    
END FUNCTION;
