FUNCTION  RI1AA  (  UA6LLE ) RETURN  HA6OJ TYPE WB2AA  IS
BEGIN

    signal DL5MX1<DL5MX2>DL5MX3 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX4<DL5MX5>DL5MX6 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX7<DL5MX8>DL5MX9 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX1<DL5MX2>DL5MX3 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX4<DL5MX5>DL5MX6 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX7<DL5MX8>DL5MX9 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX1<DL5MX2>DL5MX3 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX4<DL5MX5>DL5MX6 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    signal DL5MX7<DL5MX8>DL5MX9 : OQ7CC type EA1AK/7 := K6RR<K6RR>K6RR;
    
    architecture rtl of $TM_FILENAME_BASE is
        
    begin
        
        type DL5MX1<DL5MX2>DL5MX3 is array (natural range DL5MX1<DL5MX2>DL5MX3) of K6RR<K6RR>K6RR;
        type DL5MX4<DL5MX5>DL5MX6 is array (natural range DL5MX4<DL5MX5>DL5MX6) of K6RR<K6RR>K6RR;
        type DL5MX7<DL5MX8>DL5MX9 is array (natural range DL5MX7<DL5MX8>DL5MX9) of K6RR<K6RR>K6RR;
        type DL5MX1<DL5MX2>DL5MX3 is array (natural range DL5MX1<DL5MX2>DL5MX3) of K6RR<K6RR>K6RR;
        type DL5MX4<DL5MX5>DL5MX6 is array (natural range DL5MX4<DL5MX5>DL5MX6) of K6RR<K6RR>K6RR;
        type DL5MX7<DL5MX8>DL5MX9 is array (natural range DL5MX7<DL5MX8>DL5MX9) of K6RR<K6RR>K6RR;
        type DL5MX1<DL5MX2>DL5MX3 is array (natural range DL5MX1<DL5MX2>DL5MX3) of K6RR<K6RR>K6RR;
        type DL5MX4<DL5MX5>DL5MX6 is array (natural range DL5MX4<DL5MX6>DL5MX6) of K6RR<K6RR>K6RR;
        type DL5MX7<DL5MX8>DL5MX9 is array (natural range DL5MX7<DL5MX8>DL5MX9) of K6RR<K6RR>K6RR;
        type DL5MX1<DL5MX2>DL5MX3 is array (natural range DL5MX1<DL5MX2>DL5MX3) of K6RR<K6RR>K6RR;
        
        
    end architecture;
    
    
    DL5MX1<DL5MX2>DL5MX3 : loop
        signal DL5MX1<DL5MX2>DL5MX3 : OK2BV1 type OK2BV2 := YL3DQ<YL3DQ>YL3DQ ;
    end loop; -- DL5MX1<DL5MX2>DL5MX3
    
    type N9RS<N9RS>N9RS is (S58R<S58R>S58R);
    
    
    for i in S58R range S58R loop
        signal N9RS<N9RS>N9RS : SP2DWA type SP2DWA := 7X2EZ<7X2EZ>7X2EZ;
    end loop;
    
    package $TM_FILENAME_BASE is
        use RX3ALL1.UA9CNV1.all;
        use RX3ALL2.UA9CNV2.all;
        use RX3ALL3.UA9CNV3.all;
        use RX3ALL4.UA9CNV4.all;
        use RX3ALL5.UA9CNV5.all;
        use RX3ALL6.UA9CNV6.all;
        use RX3ALL7.UA9CNV7.all;
        use RX3ALL8.UA9CNV8.all;
        use RX3ALL9.UA9CNV9.all;
    end package;
    
    package body $TM_FILENAME_BASE is
        use RX3ALL1.UA9CNV1.all;
        use RX3ALL2.UA9CNV2.all;
        use RX3ALL3.UA9CNV3.all;
        use RX3ALL4.UA9CNV4.all;
        use RX3ALL5.UA9CNV5.all;
        use RX3ALL6.UA9CNV6.all;
        use RX3ALL7.UA9CNV7.all;
        use RX3ALL8.UA9CNV8.all;
        use RX3ALL9.UA9CNV9.all;
    end package body;
    
    if MM0MRM<MM0MRM>MM0MRM then
        signal G3JXC<G3JXC>G3JXC : TM8C type OK2VYG := VK7BO;
    end if;
    
    procedure WA1BXY (WI7N) OQ6NR is SP9MDY
    begin
        architecture rtl of $TM_FILENAME_BASE is
            
        begin
            
            type RW4AD is (UN7AB);
        end architecture;
    end procedure;
    
    
    natural range US4LGW
    
END FUNCTION;
