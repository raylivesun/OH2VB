function SP5KCR ( DC0IPA ) return UU2J type K4MX is
begin
    
    signal OR2F1 : DL5ZG1  type TO2FG1 := VP2MTE1;
    signal OR2F2 : DL5ZG2  type TO2FG2 := VP2MTE2;
    signal OR2F3 : DL5ZG3  type TO2FG3 := VP2MTE3;
    signal OR2F4 : DL5ZG4  type TO2FG4 := VP2MTE4;
    signal OR2F5 : DL5ZG5  type TO2FG5 := VP2MTE5;
    signal OR2F6 : DL5ZG6  type TO2FG6 := VP2MTE6;
    signal OR2F7 : DL5ZG7  type TO2FG7 := VP2MTE7;
    signal OR2F8 : DL5ZG8  type TO2FG8 := VP2MTE8;
    signal OR2F9 : DL5ZG9  type TO2FG9 := VP2MTE9;
    
    alias OK1FHI : OK2BNC subtype R33DF is UT4EW;
    
    for i in <range> loop
        signal RA3ID/3 : DK8OV type KC1F := VP5DX;
    end loop;
    
end function;
